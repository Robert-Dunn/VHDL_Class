library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE ieee.numeric_std.ALL;

entity digital_to_distance is
Port(
	clk : in STD_LOGIC;
	reset: in STD_LOGIC;
	done: in STD_LOGIC;
	binary_input: in STD_LOGIC_VECTOR (7 downto 0);
	switches: in STD_LOGIC_VECTOR(1 downto 0);
	tens: out integer;
	ones: out integer;
	tenths: out integer;
	hundredths: out integer
);
end digital_to_distance;

architecture Behavioral of digital_to_distance is

type digits is array (0 to 170,1 to 8)of integer;
constant LUT: digits := --first four digits is cm next four inches 
((3,0,0,9,1,1,8,5),
(2,9,2,8,1,1,5,3),
(2,8,5,0,1,1,2,2),
(2,7,7,5,1,0,9,3),
(2,7,0,4,1,0,6,4),
(2,6,3,5,1,0,3,7),
(2,5,7,0,1,0,1,2),
(2,5,0,7,0,9,8,7),
(2,4,4,6,0,9,6,3),
(2,3,8,8,0,9,4,0),
(2,3,3,3,0,9,1,9),
(2,2,8,0,0,8,9,8),
(2,2,2,9,0,8,7,8),
(2,1,8,0,0,8,5,8),
(2,1,3,3,0,8,4,0),
(2,0,8,8,0,8,2,2),
(2,0,4,5,0,8,0,5),
(2,0,0,3,0,7,8,9),
(1,9,6,3,0,7,7,3),
(1,9,2,5,0,7,5,8),
(1,8,8,8,0,7,4,3),
(1,8,5,2,0,7,2,9),
(1,8,1,8,0,7,1,6),
(1,7,8,5,0,7,0,3),
(1,7,5,3,0,6,9,0),
(1,7,2,2,0,6,7,8),
(1,6,9,3,0,6,6,6),
(1,6,6,4,0,6,5,5),
(1,6,3,7,0,6,4,4),
(1,6,1,0,0,6,3,4),
(1,5,8,4,0,6,2,4),
(1,5,5,9,0,6,1,4),
(1,5,3,5,0,6,0,4),
(1,5,1,1,0,5,9,5),
(1,4,8,8,0,5,8,6),
(1,4,6,6,0,5,7,7),
(1,4,4,5,0,5,6,9),
(1,4,2,4,0,5,6,1),
(1,4,0,4,0,5,5,3),
(1,3,8,4,0,5,4,5),
(1,3,6,4,0,5,3,7),
(1,3,4,6,0,5,3,0),
(1,3,2,7,0,5,2,3),
(1,3,0,9,0,5,1,6),
(1,2,9,2,0,5,0,9),
(1,2,7,5,0,5,0,2),
(1,2,5,8,0,4,9,5),
(1,2,4,2,0,4,8,9),
(1,2,2,6,0,4,8,3),
(1,2,1,0,0,4,7,6),
(1,1,9,5,0,4,7,0),
(1,1,8,0,0,4,6,4),
(1,1,6,5,0,4,5,9),
(1,1,5,1,0,4,5,3),
(1,1,3,6,0,4,4,7),
(1,1,2,2,0,4,4,2),
(1,1,0,9,0,4,3,7),
(1,0,9,5,0,4,3,1),
(1,0,8,2,0,4,2,6),
(1,0,6,9,0,4,2,1),
(1,0,5,7,0,4,1,6),
(1,0,4,4,0,4,1,1),
(1,0,3,2,0,4,0,6),
(1,0,2,0,0,4,0,2),
(1,0,0,8,0,3,9,7),
(0,9,9,7,0,3,9,2),
(0,9,8,5,0,3,8,8),
(0,9,7,4,0,3,8,3),
(0,9,6,3,0,3,7,9),
(0,9,5,2,0,3,7,5),
(0,9,4,2,0,3,7,1),
(0,9,3,1,0,3,6,7),
(0,9,2,1,0,3,6,3),
(0,9,1,1,0,3,5,9),
(0,9,0,2,0,3,5,5),
(0,8,9,2,0,3,5,1),
(0,8,8,3,0,3,4,7),
(0,8,7,3,0,3,4,4),
(0,8,6,4,0,3,4,0),
(0,8,5,6,0,3,3,7),
(0,8,4,7,0,3,3,3),
(0,8,3,9,0,3,3,0),
(0,8,3,0,0,3,2,7),
(0,8,2,2,0,3,2,4),
(0,8,1,5,0,3,2,1),
(0,8,0,7,0,3,1,8),
(0,7,9,9,0,3,1,5),
(0,7,9,2,0,3,1,2),
(0,7,8,5,0,3,0,9),
(0,7,7,8,0,3,0,6),
(0,7,7,1,0,3,0,4),
(0,7,6,5,0,3,0,1),
(0,7,5,8,0,2,9,9),
(0,7,5,2,0,2,9,6),
(0,7,4,6,0,2,9,4),
(0,7,4,0,0,2,9,1),
(0,7,3,4,0,2,8,9),
(0,7,2,9,0,2,8,7),
(0,7,2,3,0,2,8,5),
(0,7,1,8,0,2,8,3),
(0,7,1,3,0,2,8,1),
(0,7,0,7,0,2,7,9),
(0,7,0,2,0,2,7,7),
(0,6,9,8,0,2,7,5),
(0,6,9,3,0,2,7,3),
(0,6,8,8,0,2,7,1),
(0,6,8,4,0,2,6,9),
(0,6,7,9,0,2,6,7),
(0,6,7,5,0,2,6,6),
(0,6,7,1,0,2,6,4),
(0,6,6,6,0,2,6,2),
(0,6,6,2,0,2,6,1),
(0,6,5,8,0,2,5,9),
(0,6,5,4,0,2,5,8),
(0,6,5,0,0,2,5,6),
(0,6,4,6,0,2,5,4),
(0,6,4,2,0,2,5,3),
(0,6,3,9,0,2,5,1),
(0,6,3,5,0,2,5,0),
(0,6,3,1,0,2,4,8),
(0,6,2,7,0,2,4,7),
(0,6,2,3,0,2,4,5),
(0,6,1,9,0,2,4,4),
(0,6,1,5,0,2,4,2),
(0,6,1,1,0,2,4,1),
(0,6,0,7,0,2,3,9),
(0,6,0,3,0,2,3,8),
(0,5,9,9,0,2,3,6),
(0,5,9,5,0,2,3,4),
(0,5,9,1,0,2,3,3),
(0,5,8,7,0,2,3,1),
(0,5,8,2,0,2,2,9),
(0,5,7,8,0,2,2,8),
(0,5,7,4,0,2,2,6),
(0,5,6,9,0,2,2,4),
(0,5,6,4,0,2,2,2),
(0,5,6,0,0,2,2,0),
(0,5,5,5,0,2,1,8),
(0,5,5,0,0,2,1,7),
(0,5,4,5,0,2,1,5),
(0,5,4,0,0,2,1,3),
(0,5,3,5,0,2,1,1),
(0,5,3,0,0,2,0,8),
(0,5,2,4,0,2,0,6),
(0,5,1,9,0,2,0,4),
(0,5,1,3,0,2,0,2),
(0,5,0,8,0,2,0,0),
(0,5,0,2,0,1,9,8),
(0,4,9,7,0,1,9,6),
(0,4,9,1,0,1,9,3),
(0,4,8,5,0,1,9,1),
(0,4,8,0,0,1,8,9),
(0,4,7,4,0,1,8,7),
(0,4,6,8,0,1,8,4),
(0,4,6,3,0,1,8,2),
(0,4,5,7,0,1,8,0),
(0,4,5,1,0,1,7,8),
(0,4,4,6,0,1,7,6),
(0,4,4,1,0,1,7,4),
(0,4,3,6,0,1,7,2),
(0,4,3,1,0,1,7,0),
(0,4,2,6,0,1,6,8),
(0,4,2,2,0,1,6,6),
(0,4,1,7,0,1,6,4),
(0,4,1,4,0,1,6,3),
(0,4,1,0,0,1,6,1),
(0,4,0,7,0,1,6,0),
(0,4,0,4,0,1,5,9),
(0,4,0,2,0,1,5,8),
(0,4,0,1,0,1,5,8),
(0,4,0,0,0,1,5,7));

signal integer_input: integer;

begin

Distance : process(clk,switches,reset)
variable index: integer;
variable ten: integer;
variable one: integer;
variable tenth: integer;
variable hundredth: integer;
begin
	if (reset ='1') then
		ten := 0;
		one := 0;
		tenth := 0;
		hundredth := 0;	
	elsif(done = '1') then
	integer_input<=to_integer(unsigned(binary_input));
		if(integer_input >= 34 and integer_input <= 204) then
		index:=(integer_input-34);
			if(switches <="10")then 
				ten:= LUT(index,1);
				one:=LUT(index,2);
				tenth:=LUT(index,3);
				hundredth:=LUT(index,4);
			elsif(switches = "11")	then
				ten:=LUT(index,5);
				one:=LUT(index,6);
				tenth:=LUT(index,7);
				hundredth:=LUT(index,8);	
			end if;
		elsif(integer_input < 34) then
		index:= 0;
			if(switches <="10")then 
				ten:=LUT(index,1);
				one:=LUT(index,2);
				tenth:=LUT(index,3);
				hundredth:=LUT(index,4);		
			elsif(switches = "11")	then
				ten:=LUT(index,5);
				one:=LUT(index,6);
				tenth:=LUT(index,7);
				hundredth:=LUT(index,8);	
			end if;
		elsif(integer_input > 204) then
		index:= 170;
			if(switches <="10")then 
				ten:=LUT(index,1);
				one:=LUT(index,2);
				tenth:=LUT(index,3);
				hundredth:=LUT(index,4);
			elsif(switches = "11")	then
				ten:=LUT(index,5);
				one:=LUT(index,6);
				tenth:=LUT(index,7);
				hundredth:=LUT(index,8);			
			end if;
		end if;
	end if;
	tens <= ten;
	ones <= one;
	tenths <= tenth;
	hundredths <= hundredth;
end process;	
end Behavioral;





